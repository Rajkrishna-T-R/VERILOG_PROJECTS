`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Rajkrishna T R, Neha Fathima S
// 
// Create Date: 22.07.2025 21:10:41
// Design Name: 
// Module Name: mod_10_counter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: Counter which can count till  a certain number (here 0-9) in synchronism with one clock signal,
//              It has a set time mode which will hold the count 
//              During set time mode if select (slt) signal is activated, it will count with in synchronism with another clock signal  
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mod_10_counter(

                      count,
                      
                      carry,
                      
                      clear,
                      
                      clkmain,
                      
                      slt,
                      
                      set_time
                      
                      
                      );



input clkmain;    // Main clock T = 1s

input slt;     // for selectively accessing this counter

input set_time;   // for time setting

input clear;      // for clearing count

output reg [3:0]count; // count 4 bit 

output reg carry;      // carry for subsequent digit

always@(posedge clkmain  or posedge clear)
 
 begin
 
    if(clear==1'b1)     // major condition
      
      begin 
      
        count<=4'd0;
        
        carry<=1'b0;
      
      end
        
      else if (set_time == 1'b1 && slt == 1'b0)
      
       begin
             // Hold mode 
             
             count <= count;  
             
             carry <= 1'b0;
             
       end     
       
      else if(slt>1'b0 && set_time>1'b0) // time setting mode
       
        begin
            
           if(count>=4'd9)   // counting for setting time
           
               begin
            
                count<=4'd0;
                
                carry<=1'b1;
               
               end
            
           else 
            
                begin
                    
                    count<=count+1'b1;  //counting for setting time
                    
                    carry<=1'b0;
                    
                end
            
        end   
        
     else if (count>=4'd9)          // normal carry 
            
            begin
                     
                count<=4'd0;
                
                carry<=1'b1;
        
            end
        
     else                             // Normal operation 
            
            begin
                
                count<=count+1'b1;
                
                carry<=1'b0;
                
                
            end
    end
  
endmodule